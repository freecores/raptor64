module Raptor64_tb();
parameter IDLE = 8'd1;
parameter DOCMD = 8'd2;

reg clk;
reg rst;
reg nmi;
wire sys_cyc;
wire sys_stb;
wire sys_we;
wire [7:0] sys_sel;
wire [63:0] sys_adr;
wire [63:0] sys_dbo;
wire [63:0] sys_dbi;
wire sys_ack;
reg [7:0] cnt;
wire wr_empty = 1'b1;
wire wr_full;
reg [63:0] romout;
wire stk_ack;
wire scr_ack;
wire [63:0] stk_dato;
wire [63:0] scr_dato;
wire [15:0] tc_dato;
wire tc_ack;

assign sys_ack = sys_stb|stk_ack|scr_ack|tc_ack;

initial begin
	clk = 1;
	rst = 0;
	nmi = 0;
	#100 rst = 1;
	#100 rst = 0;
	#800 nmi = 1;
	#100 nmi = 0;
end

always #10 clk = ~clk;	//  50 MHz

rtfTextController tc1
(
	.rst_i(rst),
	.clk_i(clk),
	.cyc_i(sys_cyc),
	.stb_i(sys_stb),
	.ack_o(tc_ack),
	.we_i(sys_we),
	.sel_i(sys_sel[1:0]|sys_sel[3:2]|sys_sel[5:4]|sys_sel[7:6]),
	.adr_i(sys_adr),
	.dat_i(sys_dbo[15:0]),
	.dat_o(tc_dato),
	.lp(),
	.curpos(),
	.vclk(),
	.eol(),
	.eof(),
	.blank(),
	.border(),
	.rgbIn(),
	.rgbOut()
);

scratchmem u_sc
(
	.clk_i(clk),
	.cyc_i(sys_cyc),
	.stb_i(sys_stb),
	.ack_o(scr_ack),
	.we_i(sys_we),
	.sel_i(sys_sel),
	.adr_i(sys_adr),
	.dat_i(sys_dbo),
	.dat_o(scr_dato)
);

stkmem u_stk
(
	.clk_i(clk),
	.cyc_i(sys_cyc),
	.stb_i(sys_stb),
	.ack_o(stk_ack),
	.we_i(sys_we),
	.adr_i(sys_adr),
	.dat_i(sys_dbo),
	.dat_o(stk_dato)
);

reg [63:0] keybdout;
always @(sys_adr)
	if (sys_adr==64'hFFFF_FFFF_FFDC_0000) begin
		$display ("keyboard=FF");
		keybdout <= 64'hFFFF_FFFF_FFFF_FFFF;
	end
	else
		keybdout <= 64'd0;
	
always @(sys_adr)
case(sys_adr)// | 64'hFFFF_FFFF_FFFF_0000)
64'hFFFFFFFFFFFFF000:	romout <= 64'h000030000000000A;
64'hFFFFFFFFFFFFF008:	romout <= 64'h0BEFFFFEFF800000;
64'hFFFFFFFFFFFFF010:	romout <= 64'h001050A3000000CE;
64'hFFFFFFFFFFFFF018:	romout <= 64'h1080600041462018;
64'hFFFFFFFFFFFFF020:	romout <= 64'h001058A300000020;
64'hFFFFFFFFFFFFF028:	romout <= 64'h1080400041662018;
64'hFFFFFFFFFFFFF030:	romout <= 64'h000036F886000048;
64'hFFFFFFFFFFFFF038:	romout <= 64'h1080600041400000;
64'hFFFFFFFFFFFFF040:	romout <= 64'h001060C7FFFFFCC6;
64'hFFFFFFFFFFFFF048:	romout <= 64'h1880000041A62000;
64'hFFFFFFFFFFFFF050:	romout <= 64'h001070A100000001;
64'hFFFFFFFFFFFFF058:	romout <= 64'h0A1FFFFF0E060008;
64'hFFFFFFFFFFFFF060:	romout <= 64'h002AA0C7FFFFFDC1;
64'hFFFFFFFFFFFFF068:	romout <= 64'h2F84000018902008;
64'hFFFFFFFFFFFFF070:	romout <= 64'h0022A4A176543210;
64'hFFFFFFFFFFFFF078:	romout <= 64'h008400009A902100;
64'hFFFFFFFFFFFFF080:	romout <= 64'h0024A4A1FEDCBA98;
64'hFFFFFFFFFFFFF088:	romout <= 64'h00840000A2902100;
64'hFFFFFFFFFFFFF090:	romout <= 64'h000028CFFFFFFE6A;
64'hFFFFFFFFFFFFF098:	romout <= 64'h03FBC000018BE000;
64'hFFFFFFFFFFFFF0A0:	romout <= 64'hFFC3427F40000003;
64'hFFFFFFFFFFFFF0A8:	romout <= 64'h1008200000028BFF;
64'hFFFFFFFFFFFFF0B0:	romout <= 64'hFFF132F8400000A8;
64'hFFFFFFFFFFFFF0B8:	romout <= 64'h0288400000131FFF;
64'hFFFFFFFFFFFFF0C0:	romout <= 64'h00000EF801FFFF4A;
64'hFFFFFFFFFFFFF0C8:	romout <= 64'h0DFBFE000039DD00;
64'hFFFFFFFFFFFFF0D0:	romout <= 64'h6F57206F6C6C6548;
64'hFFFFFFFFFFFFF0E0:	romout <= 64'h3436726F74706152;
64'hFFFFFFFFFFFFF0E8:	romout <= 64'h206D657473797320;
64'hFFFFFFFFFFFFF0F0:	romout <= 64'h676E697472617473;
64'hFFFFFFFFFFFFF0F8:	romout <= 64'h000000002E2E2E2E;
64'hFFFFFFFFFFFFF100:	romout <= 64'h0000003FBC000008;
64'hFFFFFFFFFFFFF108:	romout <= 64'h0A1FFDC0A0067E18;
64'hFFFFFFFFFFFFF110:	romout <= 64'h0000060046000001;
64'hFFFFFFFFFFFFF118:	romout <= 64'h2F8C000000814318;
64'hFFFFFFFFFFFFF120:	romout <= 64'h0000011F86000000;
64'hFFFFFFFFFFFFF128:	romout <= 64'h0DFBFE0000180108;
64'hFFFFFFFFFFFFF130:	romout <= 64'h0000203FBC000010;
64'hFFFFFFFFFFFFF138:	romout <= 64'h19F8600000067E10;
64'hFFFFFFFFFFFFF140:	romout <= 64'h000004A3FFDC0A00;
64'hFFFFFFFFFFFFF148:	romout <= 64'h0508400004080310;
64'hFFFFFFFFFFFFF150:	romout <= 64'h000002F881FFFFA8;
64'hFFFFFFFFFFFFF158:	romout <= 64'h11F8600000090308;
64'hFFFFFFFFFFFFF160:	romout <= 64'h8000091F84000008;
64'hFFFFFFFFFFFFF168:	romout <= 64'h03FBC00001837EFF;
64'hFFFFFFFFFFFFF170:	romout <= 64'h0011427F00000007;
64'hFFFFFFFFFFFFF178:	romout <= 64'h0504200000F42008;
64'hFFFFFFFFFFFFF180:	romout <= 64'h700000A300000440;
64'hFFFFFFFFFFFFF188:	romout <= 64'h18801DC000242017;
64'hFFFFFFFFFFFFF190:	romout <= 64'h000005A8C2200030;
64'hFFFFFFFFFFFFF198:	romout <= 64'h0504200000F08108;
64'hFFFFFFFFFFFFF1A0:	romout <= 64'h0011498802000450;
64'hFFFFFFFFFFFFF1A8:	romout <= 64'h2F84400010942010;
64'hFFFFFFFFFFFFF1B0:	romout <= 64'h00003C2084000001;
64'hFFFFFFFFFFFFF1B8:	romout <= 64'h1880400045214210;
64'hFFFFFFFFFFFFF1C0:	romout <= 64'h0000627700000007;
64'hFFFFFFFFFFFFF1C8:	romout <= 64'h000000000200BEF0;
64'hFFFFFFFFFFFFF1D0:	romout <= 64'h000001800200041C;
64'hFFFFFFFFFFFFF1D8:	romout <= 64'h03FBC000010360F8;
64'hFFFFFFFFFFFFF1E0:	romout <= 64'h7000027F40000002;
64'hFFFFFFFFFFFFF1E8:	romout <= 64'h2008200000028BFF;
64'hFFFFFFFFFFFFF1F0:	romout <= 64'h00000AF841FFFFC1;
64'hFFFFFFFFFFFFF1F8:	romout <= 64'h050420000FF80200;
64'hFFFFFFFFFFFFF200:	romout <= 64'h0002A1000400041C;
64'hFFFFFFFFFFFFF208:	romout <= 64'h2C04548000DBE200;
64'hFFFFFFFFFFFFF210:	romout <= 64'h000008C7FFFFFD2D;
64'hFFFFFFFFFFFFF218:	romout <= 64'h0DFBFE000029DD00;
64'hFFFFFFFFFFFFF220:	romout <= 64'h00000C3FBC000010;
64'hFFFFFFFFFFFFF228:	romout <= 64'h118020004009FC00;
64'hFFFFFFFFFFFFF230:	romout <= 64'h0010002042000001;
64'hFFFFFFFFFFFFF238:	romout <= 64'h0A2FFD0000066008;
64'hFFFFFFFFFFFFF240:	romout <= 64'h0000050882000066;
64'hFFFFFFFFFFFFF248:	romout <= 64'h1888200006608108;
64'hFFFFFFFFFFFFF250:	romout <= 64'h0010010801FF0000;
64'hFFFFFFFFFFFFF258:	romout <= 64'h0504200007F46008;
64'hFFFFFFFFFFFFF260:	romout <= 64'hFFF27AC840080040;
64'hFFFFFFFFFFFFF268:	romout <= 64'h2770000000331FFF;
64'hFFFFFFFFFFFFF270:	romout <= 64'h0000802FBC000010;
64'hFFFFFFFFFFFFF278:	romout <= 64'h03FBC00002000000;
64'hFFFFFFFFFFFFF280:	romout <= 64'hFFF4727F40000007;
64'hFFFFFFFFFFFFF288:	romout <= 64'h0204201000031FFF;
64'hFFFFFFFFFFFFF290:	romout <= 64'h8000110844000000;
64'hFFFFFFFFFFFFF298:	romout <= 64'h1884400000006210;
64'hFFFFFFFFFFFFF2A0:	romout <= 64'h0003211804000408;
64'hFFFFFFFFFFFFF2A8:	romout <= 64'h10806000414BE110;
64'hFFFFFFFFFFFFF2B0:	romout <= 64'h0010218886000000;
64'hFFFFFFFFFFFFF2B8:	romout <= 64'h2774000000766008;
64'hFFFFFFFFFFFFF2C0:	romout <= 64'h004FF4DFBFE00004;
64'hFFFFFFFFFFFFF2C8:	romout <= 64'h0580400042B16008;
64'hFFFFFFFFFFFFF2D0:	romout <= 64'hFFFFFC1044500018;
64'hFFFFFFFFFFFFF2D8:	romout <= 64'h05803D00000FFFFF;
64'hFFFFFFFFFFFFF2E0:	romout <= 64'h0000505804000032;
64'hFFFFFFFFFFFFF2E8:	romout <= 64'h1884400000016018;
64'hFFFFFFFFFFFFF2F0:	romout <= 64'h0000042842000002;
64'hFFFFFFFFFFFFF2F8:	romout <= 64'h2F8C1FFFFC90C318;
64'hFFFFFFFFFFFFF300:	romout <= 64'h000000C7FFFFFFFE;
64'hFFFFFFFFFFFFF308:	romout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFF310:	romout <= 64'h0000037800000000;
64'hFFFFFFFFFFFFF318:	romout <= 64'h03FBC000028DE000;
64'hFFFFFFFFFFFFF320:	romout <= 64'h6800027F4000000F;
64'hFFFFFFFFFFFFF328:	romout <= 64'h108C200000028FFF;
64'hFFFFFFFFFFFFF330:	romout <= 64'h80006108C4000002;
64'hFFFFFFFFFFFFF338:	romout <= 64'h0100440000904110;
64'hFFFFFFFFFFFFF340:	romout <= 64'hFFF430A100000020;
64'hFFFFFFFFFFFFF348:	romout <= 64'h0A3FFD0000031FFF;
64'hFFFFFFFFFFFFF350:	romout <= 64'h00000988C2000000;
64'hFFFFFFFFFFFFF358:	romout <= 64'h2F80400000F08318;
64'hFFFFFFFFFFFFF360:	romout <= 64'h0010501008200009;
64'hFFFFFFFFFFFFF368:	romout <= 64'h0A3FFD1000042008;
64'hFFFFFFFFFFFFF370:	romout <= 64'h00000988C2000000;
64'hFFFFFFFFFFFFF378:	romout <= 64'h2F80400000F08318;
64'hFFFFFFFFFFFFF380:	romout <= 64'h800016774000000F;
64'hFFFFFFFFFFFFF388:	romout <= 64'h03FBC00002837EFF;
64'hFFFFFFFFFFFFF390:	romout <= 64'h6800027F4000000F;
64'hFFFFFFFFFFFFF398:	romout <= 64'h108C200000028FFF;
64'hFFFFFFFFFFFFF3A0:	romout <= 64'h80006108C4000002;
64'hFFFFFFFFFFFFF3A8:	romout <= 64'h0108220000504110;
64'hFFFFFFFFFFFFF3B0:	romout <= 64'h000084A3FFD00000;
64'hFFFFFFFFFFFFF3B8:	romout <= 64'h188C80000006A309;
64'hFFFFFFFFFFFFF3C0:	romout <= 64'hFFFEBC28C6000002;
64'hFFFFFFFFFFFFF3C8:	romout <= 64'h0A3FFDA0000BE017;
64'hFFFFFFFFFFFFF3D0:	romout <= 64'h00000508C2000002;
64'hFFFFFFFFFFFFF3D8:	romout <= 64'h0C7FFFFFCFA0E108;
64'hFFFFFFFFFFFFF3E0:	romout <= 64'h800016774000000F;
64'hFFFFFFFFFFFFF3E8:	romout <= 64'h03FBC00001837EFF;
64'hFFFFFFFFFFFFF3F0:	romout <= 64'h6800027F00000007;
64'hFFFFFFFFFFFFF3F8:	romout <= 64'h108C400000028FFF;
64'hFFFFFFFFFFFFF400:	romout <= 64'h2000001082300018;
64'hFFFFFFFFFFFFF408:	romout <= 64'h028C7D0000006318;
64'hFFFFFFFFFFFFF410:	romout <= 64'h000000A100000020;
64'hFFFFFFFFFFFFF418:	romout <= 64'h028C600000262308;
64'hFFFFFFFFFFFFF420:	romout <= 64'h00001EF805FFFFAF;
64'hFFFFFFFFFFFFF428:	romout <= 64'h0DFBFE000039DC00;
64'hFFFFFFFFFFFFF430:	romout <= 64'h80010450420000FF;
64'hFFFFFFFFFFFFF438:	romout <= 64'h2B04020005AA8100;
64'hFFFFFFFFFFFFF440:	romout <= 64'h400186B84010007A;
64'hFFFFFFFFFFFFF448:	romout <= 64'h03042000060A8100;
64'hFFFFFFFFFFFFF450:	romout <= 64'h0000005842000100;
64'hFFFFFFFFFFFFF458:	romout <= 64'h050420000FF360F8;
64'hFFFFFFFFFFFFF460:	romout <= 64'h0000F2B84008001A;
64'hFFFFFFFFFFFFF468:	romout <= 64'h0D83E0000000A108;
64'hFFFFFFFFFFFFF470:	romout <= 64'h0001FD0802000418;
64'hFFFFFFFFFFFFF478:	romout <= 64'h0A3FFDA000014108;
64'hFFFFFFFFFFFFF480:	romout <= 64'h80006108C4000000;
64'hFFFFFFFFFFFFF488:	romout <= 64'h1080200041A04208;
64'hFFFFFFFFFFFFF490:	romout <= 64'h80000C504200007F;
64'hFFFFFFFFFFFFF498:	romout <= 64'h0188408000004208;
64'hFFFFFFFFFFFFF4A0:	romout <= 64'h40000188C4000016;
64'hFFFFFFFFFFFFF4A8:	romout <= 64'h010041000090A217;
64'hFFFFFFFFFFFFF4B0:	romout <= 64'h500034D83E000000;
64'hFFFFFFFFFFFFF4B8:	romout <= 64'h1880000041AB2100;
64'hFFFFFFFFFFFFF4C0:	romout <= 64'hD00244D83E000000;
64'hFFFFFFFFFFFFF4C8:	romout <= 64'h03FBC000008B2100;
64'hFFFFFFFFFFFFF4D0:	romout <= 64'h0010699F84000000;
64'hFFFFFFFFFFFFF4D8:	romout <= 64'h2C08018003842010;
64'hFFFFFFFFFFFFF4E0:	romout <= 64'h0010682884000001;
64'hFFFFFFFFFFFFF4E8:	romout <= 64'h11F8400000062010;
64'hFFFFFFFFFFFFF4F0:	romout <= 64'hC00240DFBFE00001;
64'hFFFFFFFFFFFFF4F8:	romout <= 64'h03FBC000008B2100;
64'hFFFFFFFFFFFFF500:	romout <= 64'h0010619F84000000;
64'hFFFFFFFFFFFFF508:	romout <= 64'h2C0BFE8000042010;
64'hFFFFFFFFFFFFF510:	romout <= 64'h0010603884000001;
64'hFFFFFFFFFFFFF518:	romout <= 64'h2F801FFFECA62010;
64'hFFFFFFFFFFFFF520:	romout <= 64'h000022C840280093;
64'hFFFFFFFFFFFFF528:	romout <= 64'h19F840000000FEF0;
64'hFFFFFFFFFFFFF530:	romout <= 64'hE00001080400041A;
64'hFFFFFFFFFFFFF538:	romout <= 64'h03884000001B02FE;
64'hFFFFFFFFFFFFF540:	romout <= 64'hFFF529880400041A;
64'hFFFFFFFFFFFFF548:	romout <= 64'h2C840340092BE007;
64'hFFFFFFFFFFFFF550:	romout <= 64'h0000003FBC000008;
64'hFFFFFFFFFFFFF558:	romout <= 64'h1080400041867E10;
64'hFFFFFFFFFFFFF560:	romout <= 64'h000006C0BF88001E;
64'hFFFFFFFFFFFFF568:	romout <= 64'h188040004180A210;
64'hFFFFFFFFFFFFF570:	romout <= 64'hD00252F801FFFBCA;
64'hFFFFFFFFFFFFF578:	romout <= 64'h03FBC000008B2100;
64'hFFFFFFFFFFFFF580:	romout <= 64'h0010699F84000000;
64'hFFFFFFFFFFFFF588:	romout <= 64'h2F8800000C842010;
64'hFFFFFFFFFFFFF590:	romout <= 64'hFFEB29880000041A;
64'hFFFFFFFFFFFFF598:	romout <= 64'h18800000418BE007;
64'hFFFFFFFFFFFFF5A0:	romout <= 64'h0000C2F801FFFA4A;
64'hFFFFFFFFFFFFF5A8:	romout <= 64'h27F4000001F0FEF0;
64'hFFFFFFFFFFFFF5B0:	romout <= 64'hFFF472C840180099;
64'hFFFFFFFFFFFFF5B8:	romout <= 64'h0100230000931FFF;
64'hFFFFFFFFFFFFF5C0:	romout <= 64'h0006A9080200041A;
64'hFFFFFFFFFFFFF5C8:	romout <= 64'h2C840680008BE000;
64'hFFFFFFFFFFFFF5D0:	romout <= 64'h0012A1080400041A;
64'hFFFFFFFFFFFFF5D8:	romout <= 64'h03884000001BE200;
64'hFFFFFFFFFFFFF5E0:	romout <= 64'hFFF471880400041A;
64'hFFFFFFFFFFFFF5E8:	romout <= 64'h0100230000931FFF;
64'hFFFFFFFFFFFFF5F0:	romout <= 64'h000009080200041A;
64'hFFFFFFFFFFFFF5F8:	romout <= 64'h188C400000042310;
64'hFFFFFFFFFFFFF600:	romout <= 64'h00000428C6000002;
64'hFFFFFFFFFFFFF608:	romout <= 64'h0A4FFDA00000A108;
64'hFFFFFFFFFFFFF610:	romout <= 64'hFFFC92090A000000;
64'hFFFFFFFFFFFFF618:	romout <= 64'h0A200000020BE12F;
64'hFFFFFFFFFFFFF620:	romout <= 64'h0008A988C5FFFFFE;
64'hFFFFFFFFFFFFF628:	romout <= 64'h2C04040000ABE000;
64'hFFFFFFFFFFFFF630:	romout <= 64'hFFF4701002400009;
64'hFFFFFFFFFFFFF638:	romout <= 64'h0100230000931FFF;
64'hFFFFFFFFFFFFF640:	romout <= 64'hFFF4301008100009;
64'hFFFFFFFFFFFFF648:	romout <= 64'h188C200000031FFF;
64'hFFFFFFFFFFFFF650:	romout <= 64'h00007CC7FFFFFD9C;
64'hFFFFFFFFFFFFF658:	romout <= 64'h0DFBFE000069DD00;
64'hFFFFFFFFFFFFF660:	romout <= 64'h00007CC7FFFFFDAC;
64'hFFFFFFFFFFFFF668:	romout <= 64'h0DFBFE000069DD00;
64'hFFFFFFFFFFFFF670:	romout <= 64'h00001C3FBC000020;
64'hFFFFFFFFFFFFF678:	romout <= 64'h0A3FFDA00009FD00;
64'hFFFFFFFFFFFFF680:	romout <= 64'h00000608C2000016;
64'hFFFFFFFFFFFFF688:	romout <= 64'h248C20000160A108;
64'hFFFFFFFFFFFFF690:	romout <= 64'h000005080200041A;
64'hFFFFFFFFFFFFF698:	romout <= 64'h1880200041A0A108;
64'hFFFFFFFFFFFFF6A0:	romout <= 64'h000B1A08C4000000;
64'hFFFFFFFFFFFFF6A8:	romout <= 64'h1880000041ABE110;
64'hFFFFFFFFFFFFF6B0:	romout <= 64'h0000050802000418;
64'hFFFFFFFFFFFFF6B8:	romout <= 64'h188020004180A108;
64'hFFFFFFFFFFFFF6C0:	romout <= 64'h000008A3FFDA0000;
64'hFFFFFFFFFFFFF6C8:	romout <= 64'h2F8440001C682310;
64'hFFFFFFFFFFFFF6D0:	romout <= 64'h0010603884000001;
64'hFFFFFFFFFFFFF6D8:	romout <= 64'h108C400000062010;
64'hFFFFFFFFFFFFF6E0:	romout <= 64'h0000581884080000;
64'hFFFFFFFFFFFFF6E8:	romout <= 64'h0104410000542308;
64'hFFFFFFFFFFFFF6F0:	romout <= 64'hFFF38988C2000016;
64'hFFFFFFFFFFFFF6F8:	romout <= 64'h2774000000731FFF;
64'hFFFFFFFFFFFFF700:	romout <= 64'h000060DFBFE00004;
64'hFFFFFFFFFFFFF708:	romout <= 64'h27F400000030DEF0;
64'hFFFFFFFFFFFFF710:	romout <= 64'h0002A12844000000;
64'hFFFFFFFFFFFFF718:	romout <= 64'h0C7FFFFFD2DBE200;
64'hFFFFFFFFFFFFF720:	romout <= 64'h00000EF801FFFF8A;
64'hFFFFFFFFFFFFF728:	romout <= 64'h0DFBFE000039DD00;
64'hFFFFFFFFFFFFF730:	romout <= 64'h0000003FBC000008;
64'hFFFFFFFFFFFFF738:	romout <= 64'h0C7FFFFFDC167EF8;
64'hFFFFFFFFFFFFF740:	romout <= 64'h0000211FBE000000;
64'hFFFFFFFFFFFFF748:	romout <= 64'h037BC0000100BEF0;
64'hFFFFFFFFFFFFF750:	romout <= 64'h0000219F82000000;
64'hFFFFFFFFFFFFF758:	romout <= 64'h0A10000000D67EF8;
64'hFFFFFFFFFFFFF760:	romout <= 64'h000028C7FFFFFD2D;
64'hFFFFFFFFFFFFF768:	romout <= 64'h0C7FFFFFD2D28400;
64'hFFFFFFFFFFFFF770:	romout <= 64'h0000211F82000000;
64'hFFFFFFFFFFFFF778:	romout <= 64'h0DFBFE0000247EF8;
64'hFFFFFFFFFFFFF780:	romout <= 64'h00002037BC000010;
64'hFFFFFFFFFFFFF788:	romout <= 64'h19F8200000067EF8;
64'hFFFFFFFFFFFFF790:	romout <= 64'h0000C0504200000F;
64'hFFFFFFFFFFFFF798:	romout <= 64'h2B04014003908108;
64'hFFFFFFFFFFFFF7A0:	romout <= 64'hFFF4B42042000007;
64'hFFFFFFFFFFFFF7A8:	romout <= 64'h11F8200000031FFF;
64'hFFFFFFFFFFFFF7B0:	romout <= 64'h8000091FBE000008;
64'hFFFFFFFFFFFFF7B8:	romout <= 64'h03FBC00001037EFF;
64'hFFFFFFFFFFFFF7C0:	romout <= 64'h8000127F40000001;
64'hFFFFFFFFFFFFF7C8:	romout <= 64'h0C7FFFFFDE006108;
64'hFFFFFFFFFFFFF7D0:	romout <= 64'hFFF7801842200002;
64'hFFFFFFFFFFFFF7D8:	romout <= 64'h2774000000131FFF;
64'hFFFFFFFFFFFFF7E0:	romout <= 64'h000060DFBFE00002;
64'hFFFFFFFFFFFFF7E8:	romout <= 64'h27F400000050FEF0;
64'hFFFFFFFFFFFFF7F0:	romout <= 64'h000008A300000007;
64'hFFFFFFFFFFFFF7F8:	romout <= 64'h0C7FFFFFDEE06109;
64'hFFFFFFFFFFFFF800:	romout <= 64'h000016F806003FCF;
64'hFFFFFFFFFFFFF808:	romout <= 64'h0DFBFE000039DD00;
64'hFFFFFFFFFFFFF810:	romout <= 64'hFFF4B4A10000003A;
64'hFFFFFFFFFFFFF818:	romout <= 64'h0108010000931FFF;
64'hFFFFFFFFFFFFF820:	romout <= 64'h00001CC7FFFFFDF9;
64'hFFFFFFFFFFFFF828:	romout <= 64'h0A10000002028C00;
64'hFFFFFFFFFFFFF830:	romout <= 64'h000000C7FFFFFD2D;
64'hFFFFFFFFFFFFF838:	romout <= 64'h0C7FFFFFDEE40208;
64'hFFFFFFFFFFFFF840:	romout <= 64'hFFFD3C2884000001;
64'hFFFFFFFFFFFFF848:	romout <= 64'h0CFFFFFFDD2BE01F;
64'hFFFFFFFFFFFFF850:	romout <= 64'h0003F03FBC000030;
64'hFFFFFFFFFFFFF858:	romout <= 64'h0A20000000A9FC00;
64'hFFFFFFFFFFFFF860:	romout <= 64'hC00070A800000013;
64'hFFFFFFFFFFFFF868:	romout <= 64'h018C7E0000004110;
64'hFFFFFFFFFFFFF870:	romout <= 64'h800004194FE00000;
64'hFFFFFFFFFFFFF878:	romout <= 64'h0110E40000906420;
64'hFFFFFFFFFFFFF880:	romout <= 64'h400024194A200001;
64'hFFFFFFFFFFFFF888:	romout <= 64'h0704200000004519;
64'hFFFFFFFFFFFFF890:	romout <= 64'h000006F811FFFEAF;
64'hFFFFFFFFFFFFF898:	romout <= 64'h0194C80000006426;
64'hFFFFFFFFFFFFF8A0:	romout <= 64'h000004110C400009;
64'hFFFFFFFFFFFFF8A8:	romout <= 64'h010081000090652E;
64'hFFFFFFFFFFFFF8B0:	romout <= 64'h0003F0100A200009;
64'hFFFFFFFFFFFFF8B8:	romout <= 64'h0DFBFE000069DC00;
64'hFFFFFFFFFFFFF8C0:	romout <= 64'h0002703FBC000020;
64'hFFFFFFFFFFFFF8C8:	romout <= 64'h0A80000000F9FC00;
64'hFFFFFFFFFFFFF8D0:	romout <= 64'h0000C0504400000F;
64'hFFFFFFFFFFFFF8D8:	romout <= 64'h01885C0000016210;
64'hFFFFFFFFFFFFF8E0:	romout <= 64'h0000001908400001;
64'hFFFFFFFFFFFFF8E8:	romout <= 64'h0110A4000090632F;
64'hFFFFFFFFFFFFF8F0:	romout <= 64'hC0002418C6400001;
64'hFFFFFFFFFFFFF8F8:	romout <= 64'h0184220000104310;
64'hFFFFFFFFFFFFF900:	romout <= 64'h400026F811FFFE8F;
64'hFFFFFFFFFFFFF908:	romout <= 64'h0100620000904020;
64'hFFFFFFFFFFFFF910:	romout <= 64'h800012770000009C;
64'hFFFFFFFFFFFFF918:	romout <= 64'h03FBC00003837EFF;
64'hFFFFFFFFFFFFF920:	romout <= 64'hC000267F400007C4;
64'hFFFFFFFFFFFFF928:	romout <= 64'h0C7FFFFFE1404012;
64'hFFFFFFFFFFFFF930:	romout <= 64'hFFF8C01004A00009;
64'hFFFFFFFFFFFFF938:	romout <= 64'h0A90000000131FFF;
64'hFFFFFFFFFFFFF940:	romout <= 64'h600000A800000007;
64'hFFFFFFFFFFFFF948:	romout <= 64'h029CE00000006938;
64'hFFFFFFFFFFFFF950:	romout <= 64'h0003FC29CE000004;
64'hFFFFFFFFFFFFF958:	romout <= 64'h1A9D630003014118;
64'hFFFFFFFFFFFFF960:	romout <= 64'hFFFCBC1842400001;
64'hFFFFFFFFFFFFF968:	romout <= 64'h01004100009BE047;
64'hFFFFFFFFFFFFF970:	romout <= 64'h400026F813FFFE8F;
64'hFFFFFFFFFFFFF978:	romout <= 64'h0C7FFFFFE3004050;
64'hFFFFFFFFFFFFF980:	romout <= 64'h0003FCA800000003;
64'hFFFFFFFFFFFFF988:	romout <= 64'h1AA1630003014118;
64'hFFFFFFFFFFFFF990:	romout <= 64'hFFFEBC1842400001;
64'hFFFFFFFFFFFFF998:	romout <= 64'h182C0000014BE047;
64'hFFFFFFFFFFFFF9A0:	romout <= 64'h80001E77400007C4;
64'hFFFFFFFFFFFFF9A8:	romout <= 64'h0C7FFFFFDD237EFF;
64'hFFFFFFFFFFFFF9B0:	romout <= 64'hFFF4B4A100000024;
64'hFFFFFFFFFFFFF9B8:	romout <= 64'h0C7FFFFFC7631FFF;
64'hFFFFFFFFFFFFF9C0:	romout <= 64'hFFF4B6C04010000D;
64'hFFFFFFFFFFFFF9C8:	romout <= 64'h2F801FFFFCA31FFF;
64'hFFFFFFFFFFFFF9D0:	romout <= 64'hFFF471880000041A;
64'hFFFFFFFFFFFFF9D8:	romout <= 64'h0104030000931FFF;
64'hFFFFFFFFFFFFF9E0:	romout <= 64'h00000908C2000000;
64'hFFFFFFFFFFFFF9E8:	romout <= 64'h0C7FFFFFD160A318;
64'hFFFFFFFFFFFFF9F0:	romout <= 64'h000002C840140024;
64'hFFFFFFFFFFFFF9F8:	romout <= 64'h028C600000242308;
64'hFFFFFFFFFFFFFA00:	romout <= 64'hC000E8C7FFFFFD16;
64'hFFFFFFFFFFFFFA08:	romout <= 64'h2C041800044B0104;
64'hFFFFFFFFFFFFFA10:	romout <= 64'h50012AC075F00042;
64'hFFFFFFFFFFFFFA18:	romout <= 64'h2C045E8004CB0105;
64'hFFFFFFFFFFFFFA20:	romout <= 64'h40010EC04044003F;
64'hFFFFFFFFFFFFFA28:	romout <= 64'h2F801FFFC4AB0100;
64'hFFFFFFFFFFFFFA30:	romout <= 64'h00000908C2000000;
64'hFFFFFFFFFFFFFA38:	romout <= 64'h0C7FFFFFD160A318;
64'hFFFFFFFFFFFFFA40:	romout <= 64'h000002C87F68004C;
64'hFFFFFFFFFFFFFA48:	romout <= 64'h028C600000242308;
64'hFFFFFFFFFFFFFA50:	romout <= 64'h60014CC7FFFFFD16;
64'hFFFFFFFFFFFFFA58:	romout <= 64'h0C7FFFFFCC6B21FD;
64'hFFFFFFFFFFFFFA60:	romout <= 64'hFFE9C2F801FFFA4A;
64'hFFFFFFFFFFFFFA68:	romout <= 64'h0C7FFFFFDC1287FF;
64'hFFFFFFFFFFFFFA70:	romout <= 64'h70736944203D203F;
64'hFFFFFFFFFFFFFA78:	romout <= 64'h706C65682079616C;
64'hFFFFFFFFFFFFFA80:	romout <= 64'h203D20534C430A0D;
64'hFFFFFFFFFFFFFA88:	romout <= 64'h6373207261656C63;
64'hFFFFFFFFFFFFFA90:	romout <= 64'h203A0A0D6E656572;
64'hFFFFFFFFFFFFFA98:	romout <= 64'h6D2074696445203D;
64'hFFFFFFFFFFFFFAA0:	romout <= 64'h79622079726F6D65;
64'hFFFFFFFFFFFFFAA8:	romout <= 64'h3D204C0A0D736574;
64'hFFFFFFFFFFFFFAB0:	romout <= 64'h31532064616F4C20;
64'hFFFFFFFFFFFFFAB8:	romout <= 64'h0A0D656C69662039;
64'hFFFFFFFFFFFFFAC0:	romout <= 64'h706D7544203D2044;
64'hFFFFFFFFFFFFFAC8:	romout <= 64'h0D79726F6D656D20;
64'hFFFFFFFFFFFFFAD0:	romout <= 64'h617473203D20420A;
64'hFFFFFFFFFFFFFAD8:	romout <= 64'h20796E6974207472;
64'hFFFFFFFFFFFFFAE0:	romout <= 64'h4A0A0D6369736162;
64'hFFFFFFFFFFFFFAE8:	romout <= 64'h20706D754A203D20;
64'hFFFFFFFFFFFFFAF0:	romout <= 64'h0D65646F63206F74;
64'hFFFFFFFFFFFFFAF8:	romout <= 64'h000000000000000A;
64'hFFFFFFFFFFFFFB00:	romout <= 64'h0000003FBC000008;
64'hFFFFFFFFFFFFFB08:	romout <= 64'h108C200000067EF8;
64'hFFFFFFFFFFFFFB10:	romout <= 64'hFFF45828C6000002;
64'hFFFFFFFFFFFFFB18:	romout <= 64'h2C07FF0002031FFF;
64'hFFFFFFFFFFFFFB20:	romout <= 64'h00000038C6000002;
64'hFFFFFFFFFFFFFB28:	romout <= 64'h0DFBFE0000147EF8;
64'hFFFFFFFFFFFFFB30:	romout <= 64'hFFFBC4C7FFFFFEC0;
64'hFFFFFFFFFFFFFB38:	romout <= 64'h0104050000931FFF;
64'hFFFFFFFFFFFFFB40:	romout <= 64'hFFFB00A400000007;
64'hFFFFFFFFFFFFFB48:	romout <= 64'h0C7FFFFFEF131FFF;
64'hFFFFFFFFFFFFFB50:	romout <= 64'h0000058142000000;
64'hFFFFFFFFFFFFFB58:	romout <= 64'h2F809FFFFAF0A528;
64'hFFFFFFFFFFFFFB60:	romout <= 64'hFFFB02F801FFF24A;
64'hFFFFFFFFFFFFFB68:	romout <= 64'h0C7FFFFFEF131FFF;
64'hFFFFFFFFFFFFFB70:	romout <= 64'h0000001040300009;
64'hFFFFFFFFFFFFFB78:	romout <= 64'h2F801FFF1CA343F8;
64'hFFFFFFFFFFFFFB80:	romout <= 64'hFFFBC4C7FFFFFEC0;
64'hFFFFFFFFFFFFFB88:	romout <= 64'h0104020000931FFF;
64'hFFFFFFFFFFFFFB90:	romout <= 64'hFFF810C7FFFFFDD2;
64'hFFFFFFFFFFFFFB98:	romout <= 64'h0C7FFFFFE0431FFF;
64'hFFFFFFFFFFFFFBA0:	romout <= 64'hFFF810C7FFFFFE04;
64'hFFFFFFFFFFFFFBA8:	romout <= 64'h0C7FFFFFE0431FFF;
64'hFFFFFFFFFFFFFBB0:	romout <= 64'hFFF810C7FFFFFE04;
64'hFFFFFFFFFFFFFBB8:	romout <= 64'h0C7FFFFFE0431FFF;
64'hFFFFFFFFFFFFFBC0:	romout <= 64'h000062F801FFEF4A;
64'hFFFFFFFFFFFFFBC8:	romout <= 64'h27F4000000A0FEF0;
64'hFFFFFFFFFFFFFBD0:	romout <= 64'h00003CA200000000;
64'hFFFFFFFFFFFFFBD8:	romout <= 64'h108C200000029000;
64'hFFFFFFFFFFFFFBE0:	romout <= 64'hFFF45828C6000002;
64'hFFFFFFFFFFFFFBE8:	romout <= 64'h0C7FFFFFF0631FFF;
64'hFFFFFFFFFFFFFBF0:	romout <= 64'h800002C0401BFFFF;
64'hFFFFFFFFFFFFFBF8:	romout <= 64'h0504200000F06210;
64'hFFFFFFFFFFFFFC00:	romout <= 64'hFFFB3C1082200009;
64'hFFFFFFFFFFFFFC08:	romout <= 64'h01080100009BE027;
64'hFFFFFFFFFFFFFC10:	romout <= 64'h80000E774000000A;
64'hFFFFFFFFFFFFFC18:	romout <= 64'h2A04054003037EFF;
64'hFFFFFFFFFFFFFC20:	romout <= 64'h0000C2B840100039;
64'hFFFFFFFFFFFFFC28:	romout <= 64'h0D83E0000000E108;
64'hFFFFFFFFFFFFFC30:	romout <= 64'h60011AA040340041;
64'hFFFFFFFFFFFFFC38:	romout <= 64'h03842000041AE100;
64'hFFFFFFFFFFFFFC40:	romout <= 64'h000000284200000A;
64'hFFFFFFFFFFFFFC48:	romout <= 64'h2A040240061360F8;
64'hFFFFFFFFFFFFFC50:	romout <= 64'h000186B840140066;
64'hFFFFFFFFFFFFFC58:	romout <= 64'h0284200000A0E108;
64'hFFFFFFFFFFFFFC60:	romout <= 64'hFFFFFCD83E000000;
64'hFFFFFFFFFFFFFC68:	romout <= 64'h0D83E000000287FF;
64'hFFFFFFFFFFFFFC70:	romout <= 64'hAAAB541000800009;
64'hFFFFFFFFFFFFFC78:	romout <= 64'h05802AA5555F5554;
64'hFFFFFFFFFFFFFC80:	romout <= 64'h0000019A02000000;
64'hFFFFFFFFFFFFFC88:	romout <= 64'h0104430000646810;
64'hFFFFFFFFFFFFFC90:	romout <= 64'h000022F8C00000A9;
64'hFFFFFFFFFFFFFC98:	romout <= 64'h042060000000A840;
64'hFFFFFFFFFFFFFCA0:	romout <= 64'h800026F8C1FFFF00;
64'hFFFFFFFFFFFFFCA8:	romout <= 64'h0100080000904802;
64'hFFFFFFFFFFFFFCB0:	romout <= 64'hA955551A04000000;
64'hFFFFFFFFFFFFFCB8:	romout <= 64'h2F8C00001091021A;
64'hFFFFFFFFFFFFFCC0:	romout <= 64'h0000002210000008;
64'hFFFFFFFFFFFFFCC8:	romout <= 64'h2F8C1FFFF801081C;
64'hFFFFFFFFFFFFFCD0:	romout <= 64'h000026FA14000329;
64'hFFFFFFFFFFFFFCD8:	romout <= 64'h3AAAAD5552A04002;
64'hFFFFFFFFFFFFFCE0:	romout <= 64'h000000580355AAAA;
64'hFFFFFFFFFFFFFCE8:	romout <= 64'h11A0400000066808;
64'hFFFFFFFFFFFFFCF0:	romout <= 64'h0003241044300006;
64'hFFFFFFFFFFFFFCF8:	romout <= 64'h02210000008BE300;
64'hFFFFFFFFFFFFFD00:	romout <= 64'hFFFC804207000000;
64'hFFFFFFFFFFFFFD08:	romout <= 64'h01200B00009BE307;
64'hFFFFFFFFFFFFFD10:	romout <= 64'h0000001000800009;
64'hFFFFFFFFFFFFFD18:	romout <= 64'h0408755AAAA46810;
64'hFFFFFFFFFFFFFD20:	romout <= 64'h000022F8C00000A9;
64'hFFFFFFFFFFFFFD28:	romout <= 64'h0420700000008840;
64'hFFFFFFFFFFFFFD30:	romout <= 64'h000222F8C1FFFF20;
64'hFFFFFFFFFFFFFD38:	romout <= 64'h01216800014BE858;
64'hFFFFFFFFFFFFFD40:	romout <= 64'h000052FA14000048;
64'hFFFFFFFFFFFFFD48:	romout <= 64'h1981000040004852;
64'hFFFFFFFFFFFFFD50:	romout <= 64'h000080D83E000000;
64'hFFFFFFFFFFFFFD58:	romout <= 64'h0000000002000000;
64'hFFFFFFFFFFFFFD60:	romout <= 64'hFC00219803FF0000;
64'hFFFFFFFFFFFFFD68:	romout <= 64'h0080200003466017;
64'hFFFFFFFFFFFFFD70:	romout <= 64'h0008A2F841FFFFC9;
64'hFFFFFFFFFFFFFD78:	romout <= 64'h0080400042802008;
64'hFFFFFFFFFFFFFD80:	romout <= 64'hA0000408800005A9;
64'hFFFFFFFFFFFFFD88:	romout <= 64'h0104410000306211;
64'hFFFFFFFFFFFFFD90:	romout <= 64'h8000211844000000;
64'hFFFFFFFFFFFFFD98:	romout <= 64'h00880000528FFFF8;
64'hFFFFFFFFFFFFFDA0:	romout <= 64'h8000211844000008;
64'hFFFFFFFFFFFFFDA8:	romout <= 64'h008800005A8FFFF8;
64'hFFFFFFFFFFFFFDB0:	romout <= 64'h0000D40800000034;
64'hFFFFFFFFFFFFFDB8:	romout <= 64'h11803FF000002000;
64'hFFFFFFFFFFFFFDC0:	romout <= 64'h0000811805FF0008;
64'hFFFFFFFFFFFFFDC8:	romout <= 64'h3780000000000000;
64'hFFFFFFFFFFFFFFB0:	romout <= 64'h000000CFFFFFFF58;
64'hFFFFFFFFFFFFFFB8:	romout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFFFC0:	romout <= 64'h000000CFFFFFFF58;
64'hFFFFFFFFFFFFFFC8:	romout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFFFD0:	romout <= 64'h000000CFFFFFFF55;
64'hFFFFFFFFFFFFFFD8:	romout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFFFE0:	romout <= 64'h000000CFFFFFFF56;
64'hFFFFFFFFFFFFFFE8:	romout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFFFF0:	romout <= 64'h000000CFFFFFFC00;
64'hFFFFFFFFFFFFFFF8:	romout <= 64'h37800000000DE000;
default:	romout <= 64'd0;
endcase
assign sys_dbi = romout|keybdout|stk_dato|scr_dato| {4{tc_dato}};


Raptor64sc u1
(
	.rst_i(rst),
	.clk_i(clk),
	.nmi_i(nmi),
	.irq_i(1'b0),
	.bte_o(),
	.cti_o(),
	.cyc_o(sys_cyc),
	.stb_o(sys_stb),
	.ack_i(sys_ack),
	.we_o(sys_we),
	.sel_o(sys_sel),
	.adr_o(sys_adr),
	.dat_i(sys_dbi),
	.dat_o(sys_dbo),

	.sys_adv(1'b0),
	.sys_adr(59'd0)
);
endmodule
