module Raptor64_tb();
parameter IDLE = 8'd1;
parameter DOCMD = 8'd2;

reg clk;
reg rst;
reg nmi;
wire sys_cyc;
wire sys_stb;
wire sys_we;
wire [7:0] sys_sel;
wire [63:0] sys_adr;
wire [63:0] sys_dbo;
wire [63:0] sys_dbi;
wire sys_ack;
reg [7:0] cnt;
wire wr_empty = 1'b1;
wire wr_full;
reg [63:0] iromout;

assign sys_ack = sys_stb;

initial begin
	clk = 1;
	rst = 0;
	nmi = 0;
	#100 rst = 1;
	#100 rst = 0;
	#1300 nmi = 1;
	#100 nmi = 0;
end

always #10 clk = ~clk;	//  50 MHz

always @(sys_adr)
case(sys_adr)// | 64'hFFFF_FFFF_FFFF_0000)
64'hFFFFFFFFFFFFF000:	iromout <= 64'h00001CA1FFD00000;
64'hFFFFFFFFFFFFF008:	iromout <= 64'h0A30000002028800;
64'hFFFFFFFFFFFFF010:	iromout <= 64'h0000099046000000;
64'hFFFFFFFFFFFFF018:	iromout <= 64'h038840000010A108;
64'hFFFFFFFFFFFFF020:	iromout <= 64'h002AA2F881FFFF89;
64'hFFFFFFFFFFFFF028:	iromout <= 64'h2F8400001A902008;
64'hFFFFFFFFFFFFF030:	iromout <= 64'h0022A4A176543210;
64'hFFFFFFFFFFFFF038:	iromout <= 64'h008400009A902100;
64'hFFFFFFFFFFFFF040:	iromout <= 64'h0024A4A1FEDCBA98;
64'hFFFFFFFFFFFFF048:	iromout <= 64'h00840000A2902100;
64'hFFFFFFFFFFFFF050:	iromout <= 64'h004FF6F800000028;
64'hFFFFFFFFFFFFF058:	iromout <= 64'h0580400042B16008;
64'hFFFFFFFFFFFFF060:	iromout <= 64'hFFFFFC1044500018;
64'hFFFFFFFFFFFFF068:	iromout <= 64'h05803D00000FFFFF;
64'hFFFFFFFFFFFFF070:	iromout <= 64'h0000505804000032;
64'hFFFFFFFFFFFFF078:	iromout <= 64'h1884400000016018;
64'hFFFFFFFFFFFFF080:	iromout <= 64'h0000042842000002;
64'hFFFFFFFFFFFFF088:	iromout <= 64'h2F8C1FFFFC90C318;
64'hFFFFFFFFFFFFF090:	iromout <= 64'h000000C7FFFFFC2C;
64'hFFFFFFFFFFFFF098:	iromout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFF0B0:	iromout <= 64'h700003FFFFFFFFFF;
64'hFFFFFFFFFFFFF0B8:	iromout <= 64'h100440000001600F;
64'hFFFFFFFFFFFFF0C0:	iromout <= 64'h000006F881FFFFC1;
64'hFFFFFFFFFFFFF0C8:	iromout <= 64'h0D83E00000040100;
64'hFFFFFFFFFFFFF0D0:	iromout <= 64'hAAAB541000800009;
64'hFFFFFFFFFFFFF0D8:	iromout <= 64'h05802AA5555F5554;
64'hFFFFFFFFFFFFF0E0:	iromout <= 64'h0000019A02000000;
64'hFFFFFFFFFFFFF0E8:	iromout <= 64'h0104430000646810;
64'hFFFFFFFFFFFFF0F0:	iromout <= 64'h000022F8C00000A9;
64'hFFFFFFFFFFFFF0F8:	iromout <= 64'h042060000000A840;
64'hFFFFFFFFFFFFF100:	iromout <= 64'h800026F8C1FFFF00;
64'hFFFFFFFFFFFFF108:	iromout <= 64'h0100080000904802;
64'hFFFFFFFFFFFFF110:	iromout <= 64'hA955551A04000000;
64'hFFFFFFFFFFFFF118:	iromout <= 64'h2F8C00001091021A;
64'hFFFFFFFFFFFFF120:	iromout <= 64'h0000002210000008;
64'hFFFFFFFFFFFFF128:	iromout <= 64'h2F8C1FFFF801081C;
64'hFFFFFFFFFFFFF130:	iromout <= 64'h000026FA14000329;
64'hFFFFFFFFFFFFF138:	iromout <= 64'h3AAAAD5552A04002;
64'hFFFFFFFFFFFFF140:	iromout <= 64'h000000580355AAAA;
64'hFFFFFFFFFFFFF148:	iromout <= 64'h11A0400000066808;
64'hFFFFFFFFFFFFF150:	iromout <= 64'h0003241044300006;
64'hFFFFFFFFFFFFF158:	iromout <= 64'h02210000008BE300;
64'hFFFFFFFFFFFFF160:	iromout <= 64'hFFFC804207000000;
64'hFFFFFFFFFFFFF168:	iromout <= 64'h01200B00009BE307;
64'hFFFFFFFFFFFFF170:	iromout <= 64'h0000001000800009;
64'hFFFFFFFFFFFFF178:	iromout <= 64'h0408755AAAA46810;
64'hFFFFFFFFFFFFF180:	iromout <= 64'h000022F8C00000A9;
64'hFFFFFFFFFFFFF188:	iromout <= 64'h0420700000008840;
64'hFFFFFFFFFFFFF190:	iromout <= 64'h000222F8C1FFFF20;
64'hFFFFFFFFFFFFF198:	iromout <= 64'h01216800014BE858;
64'hFFFFFFFFFFFFF1A0:	iromout <= 64'h000052FA14000048;
64'hFFFFFFFFFFFFF1A8:	iromout <= 64'h1981000040004852;
64'hFFFFFFFFFFFFF1B0:	iromout <= 64'h000080D83E000000;
64'hFFFFFFFFFFFFF1B8:	iromout <= 64'h19803FF000000000;
64'hFFFFFFFFFFFFF1C0:	iromout <= 64'h0000D19805FF0008;
64'hFFFFFFFFFFFFF1C8:	iromout <= 64'h2F84000002902008;
64'hFFFFFFFFFFFFF1D0:	iromout <= 64'h0010A00802000228;
64'hFFFFFFFFFFFFF1D8:	iromout <= 64'h008800005A902010;
64'hFFFFFFFFFFFFF1E0:	iromout <= 64'h40000C1884680001;
64'hFFFFFFFFFFFFF1E8:	iromout <= 64'h1184400000004110;
64'hFFFFFFFFFFFFF1F0:	iromout <= 64'h0000200880000529;
64'hFFFFFFFFFFFFF1F8:	iromout <= 64'h008800005A946110;
64'hFFFFFFFFFFFFF200:	iromout <= 64'h0000D40800000034;
64'hFFFFFFFFFFFFF208:	iromout <= 64'h11803FF000002000;
64'hFFFFFFFFFFFFF210:	iromout <= 64'h0000811805FF0008;
64'hFFFFFFFFFFFFF218:	iromout <= 64'h3780000000000000;
64'hFFFFFFFFFFFFFFB0:	iromout <= 64'h000000CFFFFFFC6E;
64'hFFFFFFFFFFFFFFB8:	iromout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFFFC0:	iromout <= 64'h000000CFFFFFFC6E;
64'hFFFFFFFFFFFFFFC8:	iromout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFFFD0:	iromout <= 64'h0000037800000000;
64'hFFFFFFFFFFFFFFD8:	iromout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFFFE0:	iromout <= 64'h000000CFFFFFFC6D;
64'hFFFFFFFFFFFFFFE8:	iromout <= 64'h37800000000DE000;
64'hFFFFFFFFFFFFFFF0:	iromout <= 64'h000000CFFFFFFC00;
64'hFFFFFFFFFFFFFFF8:	iromout <= 64'h0000000000000000;

endcase
assign sys_dbi = iromout;


Raptor64sc u1
(
	.rst_i(rst),
	.clk_i(clk),
	.nmi_i(nmi),
	.irq_i(1'b0),
	.bte_o(),
	.cti_o(),
	.cyc_o(sys_cyc),
	.stb_o(sys_stb),
	.ack_i(sys_ack),
	.we_o(sys_we),
	.sel_o(sys_sel),
	.adr_o(sys_adr),
	.dat_i(sys_dbi),
	.dat_o(sys_dbo),

	.sys_adv(1'b0),
	.sys_adr(59'd0)
);
endmodule
